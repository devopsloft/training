#!/usr/bin/env bash

awk 'NR > 13'  README.md > challenge.md
